��n?      �sklearn.naive_bayes��MultinomialNB���)��}�(�alpha�G?�      �	fit_prior���class_prior�N�n_features_in_�M��n_features_�M��classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�class_count_�hhK ��h��R�(KK��h�f8�����R�(KhNNNJ����J����K t�b�C      *@      1@�t�b�feature_count_�hhK ��h��R�(KKM���h&�B�  �5L�4��?�����?�����W�?�m_��ǿ?�m_��ǿ?�m_��ǿ?�$Q���?9,��.��?������?qh�pZ��?�4���?����#��?�����?�����?        �W纗��?                �����?�����?��Bi���?        �V#���?�V#���?����#��?                a9c�%�?|ީ��?�����W�?�����?����#��?�����?�V#���?�����?�V#���?�����W�?�V#���?����#��?��B~�n�?        �-v�]�?        �����?��B~�n�?�����?��`�=�?����#��?�V#���?�V#���?����#��?�V#���?�m_��ǿ?�m_��ǿ?����?h��M�?        ������?�-v�]�?��B~�n�?�m_��ǿ?        �V#���?�V#���?�-v�]�?Ӈ�f�l�?�V#���?W��x��?�m_��ǿ?|�!�5�?Z���A��?�����?��`�=�?        ������?�5L�4��?WƗ�U�?        |�!�5�?�m_��ǿ?�D��	s�?��u��?�V#���?�m_��ǿ?qh�pZ��?�V#���?��eL�?                NW�FH?�?Ԕ��?����#��?�����?�����?.����?�k�=��?                �U.2]��?�V#���?�@^��V�?        7��z�?        ��`�=�?        F��d��?                        �� >� �?lx�'���?�����?N �.�?��0����?�5L�4��?�����?�V#���?�V#���?        ����?7��z�?����#��?�V#���?�V#���?        ��`�=�?        ����#��?Ѥ/�}�?                        �V#���?�����?|�!�5�?        g���>a�?        �-v�]�?B���?��`�=�?�����W�?qh�pZ��?�����?�����?        �����?�����?�����?�-v�]�?�V#���?����?�V#���?        ����#��?                �ډ��R�?        �����?������?�V#���?|�!�5�?�V#���?|�!�5�?������?7��z�?a9c�%�?�4���?��B~�n�?�4���?������?R[��N��?��z`�P�?��T	��?��$!��?        qh�pZ��?#�<����?�ER��?a9c�%�?������?�V#���?����#��?�V#���?�����?        �� >� �?        �V#���?or�N��?������?�m_��ǿ?or�N��?�V#���?        o�>����?7��z�?��`�=�?�m_��ǿ?��`�=�?�ݕd��?        ����#��?�V#���?        �����W�?        �m_��ǿ?        '�Z�p�?����#��?        �V#���?�V#���?                �V#���?7��z�?                        �V#���?��B~�n�?�m_��ǿ?                ����#��?���(,/�?�5L�4��?�*�"ps�?        c�H2g��?�����?        �4����?7��z�?        �m_��ǿ?��B~�n�?�m_��ǿ?�)�Ԁ�?�����?��B~�n�?�m_��ǿ?�V#���?��B~�n�?����#��?o�>����?�V#���?������?&�ٔ��?Ѥ/�}�?�%kS���?,���g�?qh�pZ��?��B~�n�?|�!�5�?��B~�n�?ZJ���?�m_��ǿ?        3�2�q�?�-v�]�?۪ɫ'�?�-v�]�?z���4�?�-v�]�?�����?        �����?o�>����?�$޵���?������?�$޵���?�V#���?        �4���?        �����?�V#���?�V#���?��B~�n�?�����
�?�����?                        �����W�?^i1�;�?v6{O6��?�����?�V#���?�����?�m_��ǿ?        �5L�4��?�V#���?�m_��ǿ?\���}_�? e��>*�?        \�A<��?        �m_��ǿ?�����?��T	��?�V#���?�����?�s
��?        �����?        �m_��ǿ?�m_��ǿ?�Y�O��?�����?�庖L��?        �m_����?                �����?        �����?�����?        ��`�=�?��p��?�-v�]�?        �V#���?����#��?        ������?������?�V#���?������?w5�g��?�5L�4��?        ��`�=�?�m_��ǿ?z]�4�>�?�-v�]�?        �����?�����W�?�����?���G�?�m_��ǿ?                 �-~d�?��H��?��`�=�?�m_��ǿ?        �����?�����?        ��G�a$�?'���?�V#���?�m_��ǿ?                �����?�
g�J�?�4���?����#��?����#��?�����W�?�����?��B~�n�?F��d��?7��z�?������?�����?������?�������?�m_����?�����?�4���?����#��?��f*�?�V#���?R[��N��?�V#���?�V#���?v<օ�7�?        ��p��?�bԉ�=�?�m_��ǿ?�V#���?��`�=�?����#��?�����W�?��`�=�?�:�^���?�-v�]�?                �{�M�m�?        �W纗��?�V#���?                �V#���?w5�g��?        �����?        �V#���?�m_��ǿ?�V#���?��`�=�?qh�pZ��?        pxh?�?�V#���?        ſ�a^R�?        �m_��ǿ?        |�%w�?��p��?        �����?        �s
��?        ��B~�n�?��`�=�?��Bi���?������?        �V#���?        �5L�4��?        �*+uf�?�+ ĝ�?�V#���?        �m_��ǿ?�m_��ǿ?�����
�?        0FM�G�?�����?�m_��ǿ?��ײ��?����#��?|�!�5�?�V#���?        �V#���?7��z�?�V#���?�5L�4��?�W纗��?�V#���?������?        .����?�5L�4��?�V#���?� 8֖��?�-v�]�?�m_��ǿ?�����?��`�=�?�V#���?        w5�g��?��`�=�?�5L�4��?�����?���o��?�)�I�j�?�-v�]�?|�!�5�?�m_��ǿ?�����?                                                                                                                j�"�z.�?�2�Ǔ�?�l�9Nj�?��T�?                        j�"�z.�?                        O�;�&<�?.�9�W�??���l��?                                                                                                j�"�z.�?        ǐ4۰�?                                                                                                XIVRX�?a��V��?                                O�;�&<�?                        HvE�I�?        dj)'d~@                �+p����?                r�d�O�?��s�\�?        s��,:F�? �����?                                                                �m�Z�.�?(�2W��?Gh��B�?        �/f���?                                Y�ѕ�L�?�o�����?�ἁ���?                        ����1�?         �����?        ������?        E�K���?��AnV?�?)f��?���U	�?䰉�/��?                ���N�?                                tBJ�6��?                                        [�w��%�?        {e���%�?                j�"�z.�?a��V��?rZ֞��?                        �<\L��?        E�K���?                                                        n�Wu�?                                                        �ἁ���?        bE
g�?O�;�&<�?���꼀�?{e���%�?                                                O�7�4��?        @��v���?                        m���?��?�p����?�~8����?        +>_˔�? �����?                *I�1�Q�?@��v���?                                        r�d�O�?V�Ի�?r�d�O�?        !�7�v��?��/�P��?        ���+j�?        ���y�(�?���+j�?                                        ��U�?                j�"�z.�?        tBJ�6��?        j�"�z.�?�3>`}]�?        d���?                h��=��?%_K���?                |���L�?,-�CL��?w�"��?                        ����1�?:c�}}�?                        ��8�9�?tBJ�6��?                tBJ�6��?2��EiG�?        @x,dY�?                        e�r���?                                                O�7�4��?        @��v���?                        X�DM�?                                                j�"�z.�?hG�&)�?        ��y�h��?                                �T���$�?        m���?��?                                j�"�z.�?        h��=��?                                �p����?        E�K���?��x�Z�?VF/��?                                                        tBJ�6��?                                        �<\L��?�4�.��?�a�&�z�?                                                j�"�z.�?        �<\L��?                _�y"�l @        +��Z7�?Yy6\D�?        E�K���?{e���%�?         ��r�?                O�;�&<�?        ���D�s�?        tBJ�6��?                E�K���?�^n��?                                        �<\L��?                                ��t��I�?                        ����?        tBJ�6��? �����?�Z����?�ES�w�?                w�"��?                }^�Y�?؈�����?؈�����?                <�����?��}x��?        s��,:F�?                                                                                                                                                !�7�v��?                        p�q����?@߀t��?                                                        ��Ț���?        {e���%�?�<\L��?        ʰ�aX��?g%�����?         �����?j�"�z.�?                w�"��?        �<\L��?                                        tBJ�6��?�5��?        6kC���?        tBJ�6��?        E�K���?        @߀t��?z�:��l�?        ����1�?        \��J��?                                6��H��?        �<\L��?        a��V��?�{�)���?'��"�~�?        j�"�z.�?                ��"���? �����?�Y�c���?                T��zp�?                        �<\L��?                                �2�Ǔ�?                J�4�?                        ؙ��zN�?                                        @x,dY�?                                �ꇸ�1�?��s�\�?                                �t�b�feature_log_prob_�hhK ��h��R�(KKM���h&�B�  ����������{�x����rh�����rh�����rh�����4u�%�T����WS��EvC���I����W���!�u4����"������{����{�U�"��R�S��TYp�U�"��R�U�"��R����{����{��ȉɏ�U�"��R�rZdp���$,�����"���U�"��R�U�"��R��)
k�������n�x�������{����"������{�rZdp�����{��$,��x�����$,������CX�V��0��U�"��R�a5����U�"��R����{�V��0�����{��-�ׅ�����"���h����@��$,�����"����$,��rh�����rh�����I;�s��KS	�U�"��R�EvC���a5����V��0��rh�����U�"��R��$,���$,��a5��������E���$,��C�3�o�rh�����~V{��^�ykF�������{��-�ׅ��U�"��R������������_#��U�"��R�~V{��^�rh�������k>���{�8���$,��rh�����I����W��$,��	�̂:�U�"��R�U�"��R�C�V���q�������"������{����{�'B��}���6#P��U�"��R�U�"��R��Z�rH��$,��l"_:��U�"��R��&���U�"��R��-�ׅ��U�"��R�A� j�L�U�"��R�U�"��R�U�"��R�&#3���8Q�8������{���Na��&�UY�����������{�rZdp���$,��U�"��R�I;�s��&������"���rZdp��rZdp��U�"��R��-�ׅ��U�"��R����"���֣h�;[�U�"��R�U�"��R�U�"��R��$,�����{�~V{��^�U�"��R��g�PP�U�"��R�a5����E0�J���-�ׅ���6&!5�I����W����{����{�U�"��R����{����{����{�a5�����$,��I;�s��$,��U�"��R����"���U�"��R�U�"��R��2�Ym��U�"��R����{�EvC����$,��~V{��^��$,��~V{��^�����&����)
k����!�u4�V��0����!�u4������A2�v��z�G-���g����D�I��U�"��R�I����W�N#�_L��;n����)
k��EvC����$,�����"����$,�����{�U�"��R�&#3���U�"��R��$,��N������'�ulZ�rh�����N������$,��U�"��R���u9P���&���տ{�L�rh������-�ׅ��a����5�U�"��R����"����$,��U�"��R�x����U�"��R�rh�����U�"��R�u$�[O����"���U�"��R�rZdp���$,��U�"��R�U�"��R��$,���&���U�"��R�U�"��R�U�"��R��$,��V��0��rh�����U�"��R�U�"��R����"���R!p�9��������>�gXl�U�"��R��?)+�����{�U�"��R�0� !���&���U�"��R�rh�����V��0��rh�������0n������{�V��0��rh������$,��V��0�����"�����u9P���$,�����v�����֣h�;[�L[���w,Kk?m�I����W�V��0��~V{��^�V��0��v�I�!��rh�����U�"��R��Õ(��a5�����|��a5����b�q{��a5�������{�U�"��R����{��;~���@G@E���EvC���@G@E����$,��U�"��R���!�u4�U�"��R����{��$,���$,��V��0���T�`������{�U�"��R�U�"��R�U�"��R�x������
:a��v�\0{����{��$,�����{�rh�����U�"��R���������$,��rh�������Y�7��_7[��U�"��R�'1M�B��U�"��R�rh��������{��g�����$,�����{�a�����U�"��R����{�U�"��R�rh�����rh�������*˂�����{��d�6�U�"��R���E�o�U�"��R�U�"��R����{�U�"��R����{����{�U�"��R��-�ׅ��H�s��a5����U�"��R��$,�����"���U�"��R�� Y|o���R��IV��$,���R��IV��I�&���������U�"��R��-�ׅ��rh�����%pR�36�a5����U�"��R����{�x�������{�@�x�I#�rh�����U�"��R�U�"��R�}�2r�����";��-�ׅ��rh�����U�"��R����{����{�U�"��R�������V�x)���$,��rh�����U�"��R�U�"��R����{��l������!�u4����"������"���x�������{�V��0��A� j�L��&���EvC������{�EvC����������E�o����{���!�u4����"���4�0G���$,����A2�v��$,��h����@��)2�\��U�"��R�H�s���J��yE�rh������$,���-�ׅ�����"���x�����-�ׅ���=��a5����U�"��R�U�"��R�4�5��6�U�"��R�S��TYp��$,��U�"��R�U�"��R��$,���I�&��U�"��R����{�U�"��R��$,��rh������$,���-�ׅ��I����W�U�"��R�^��[���rZdp��U�"��R������U�"��R�rh�����U�"��R���B}~�H�s��U�"��R����{�U�"��R�a�����U�"��R�V��0���-�ׅ��=���'��EvC���U�"��R��$,��U�"��R��������U�"��R�y�nS�O�|Jb�}��$,��U�"��R�rh�����rh������T�`���U�"��R�<#�V͌����{�rh�����#]N��d����"���~V{��^��$,��U�"��R��$,��ն�c��$,���������S��TYp�rZdp��EvC���U�"��R�'B��}���������$,����-b��a5����rh��������{��-�ׅ���$,��U�"��R��I�&��տ{�L�����������{�L�~��K�8�J6��a5����~V{��^�rh��������{�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�]���	���40�!u��X�b^���>��TY��{P�TY��{P�TY��{P�]���	��TY��{P�TY��{P�TY��{P��C\)Xw�����Di��֖ƈ�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�]���	��TY��{P��1k��TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P���I�w����\�		�TY��{P�TY��{P�TY��{P�TY��{P��C\)Xw�TY��{P�TY��{P�TY��{P��r��p�TY��{P����J��TY��{P�TY��{P��a��3�TY��{P�TY��{P������N�Y���=��TY��{P��'��	��:�Ra�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P��හ��b�)���� ��TY��{P�p�1�t��TY��{P�TY��{P�TY��{P�TY��{P���e�C��w�X���w�cF�TY��{P�TY��{P�TY��{P��We���TY��{P�:�Ra�TY��{P��x�����TY��{P�H�;Ň�|Ll�@n��9��k���~!��?����TY��{P�TY��{P���;�^�TY��{P�TY��{P�TY��{P�TY��{P�q����TY��{P�TY��{P�TY��{P�TY��{P�TY��{P���Kw��TY��{P��j��g]�TY��{P�TY��{P�]���	����\�		���r����TY��{P�TY��{P�TY��{P�0��s��TY��{P�H�;Ň�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P������!�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P��w�cF�TY��{P�0��m6��C\)Xw�`M�~I���j��g]�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P���)Pƌ�TY��{P�-�B�[U�TY��{P�TY��{P�TY��{P�:�o73���S<�gnJ%N��TY��{P�������:�Ra�TY��{P�TY��{P�W��-�B�[U�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P������N�Z0�c1������N�TY��{P�hC
"���X[7�TY��{P�qu�.v�TY��{P�~���5�qu�.v�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P���SI��TY��{P�TY��{P�]���	��TY��{P�q����TY��{P�]���	����q��1�TY��{P����:�:�TY��{P�TY��{P��ο��r�� ����TY��{P�TY��{P�:fa��	�D(=���\��:�TY��{P�TY��{P�TY��{P��We�������TY��{P�TY��{P�TY��{P���	���[Cs�Q%�TY��{P�TY��{P�q������{�qF�TY��{P�`�m�^�TY��{P�TY��{P�TY��{P��/WY�.�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P���)Pƌ�TY��{P�-�B�[U�TY��{P�TY��{P�TY��{P���Z�N�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�]���	���I�`��TY��{P�('VU���TY��{P�TY��{P�TY��{P�TY��{P����3H��TY��{P�:�o73��TY��{P�TY��{P�TY��{P�TY��{P�]���	��TY��{P��ο��r�TY��{P�TY��{P�TY��{P�TY��{P��S<�TY��{P�H�;Ň����v
E��.�M	�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�q����TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�0��s��ǢԖ�X�4<:�۶�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�]���	��TY��{P�0��s��TY��{P�TY��{P�Y5�ǉ��TY��{P�Z�������X��''�TY��{P�H�;Ň��j��g]�TY��{P�h��h_��TY��{P�TY��{P��C\)Xw�TY��{P����MȒ�TY��{P�q����TY��{P�TY��{P�H�;Ň��[~]�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�0��s��TY��{P�TY��{P�TY��{P�TY��{P�˗�+'��TY��{P�TY��{P�TY��{P��j-���TY��{P�q����:�Ra���]���:/,�g��TY��{P�TY��{P�\��:�TY��{P�TY��{P�D���P����gh!���gh!�TY��{P�TY��{P���ۨ���G�w�TY��{P��'��	��TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�hC
"���TY��{P�TY��{P�TY��{P�Xkl_?.�cM,v���TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P��|����TY��{P��j��g]�0��s��TY��{P��δ*�ģ��1�TY��{P�:�Ra�]���	��TY��{P�TY��{P�\��:�TY��{P�0��s��TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�q��������TY��{P���t�X�TY��{P�q����TY��{P�H�;Ň�TY��{P�cM,v������'��TY��{P��We���TY��{P��ٕh��TY��{P�TY��{P�TY��{P�TY��{P��G͎�b�TY��{P�0��s��TY��{P���\�		�qUu�[U�z]�[u��TY��{P�]���	��TY��{P�TY��{P�PK��:�Ra��R�s0�TY��{P�TY��{P���K���TY��{P�TY��{P�TY��{P�0��s��TY��{P�TY��{P�TY��{P�TY��{P�*�ؓ��TY��{P�TY��{P��2�l���TY��{P�TY��{P�TY��{P�&7�Vm�TY��{P�TY��{P�TY��{P�TY��{P�TY��{P�`�m�^�TY��{P�TY��{P�TY��{P�TY��{P�
�Xޮ��Y���=��TY��{P�TY��{P�TY��{P�TY��{P��t�b�class_log_prior_�hhK ��h��R�(KK��h&�C()i7��꿄\E��,⿔t�b�_sklearn_version��0.24.2�ub.